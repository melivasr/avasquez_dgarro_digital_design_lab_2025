module Multiplicacion32 (
    input logic [31:0] A,
    input logic [31:0] B,
    output logic [31:0] P,   // ojo: 32x32 = 64 bits
    output logic N,
    output logic Z,
    output logic C,
    output logic V
);
	logic [63:0] Pf;
	
   assign Pf = A * B;

   assign P = Pf[31:0];
	
	// Flags
   assign N = P[31];                // MSB del resultado truncado
   assign Z = (P == 32'd0);         // todo cero
   assign C = 1'b0;                 // no hay carry en mult truncada
   assign V = (Pf[63:32] != 0); // overflow si la parte alta no cabe en 32 bits
	
endmodule